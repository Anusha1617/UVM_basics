class Tx_op_mo extends uvm_monitor;


//------FACTORY Registration----------------//
	`uvm_component_utils(Tx_op_mo)

// component constructor 
function new(string name,uvm_component parent);
		super.new(name,parent);
endfunction


endclass
