gbhdff
