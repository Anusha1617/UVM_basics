mcs_dv05_ethernet_project_assertions.sv
mcs_dv05_ethernet_project_top_config.sv
mcs_dv05_ethernet_project_top.sv
